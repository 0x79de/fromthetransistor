module Processor (
    input [31:0] instruction,
    input clk,
    output [7:0] R1, R2, R3
  );
endmodule
